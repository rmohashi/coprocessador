library IEEE;
use IEEE.std_logic_1164.all;

entity reg16 is
  port (
    CLK, CLKEN, OE_L, CLR_L: in std_logic;
    D: in std_logic_vector(15 downto 0);   -- Input bus
    Q: out std_logic_vector (15 downto 0) -- Output bus (three-state)
  );
end reg16;

architecture arch of reg16 is
  signal CLR, OE: STD_LOGIC;  -- active-high versions of signals
  signal IQ: STD_LOGIC_VECTOR(15 downto 0) := (others => '0'); -- internal Q signals
begin

  process(CLK, CLR_L, CLR, OE_L, OE, IQ)
  begin
    CLR <= not CLR_L; 
	  OE <= not OE_L;

    if (CLR = '1') then
		  IQ <= (others => '0');
    elsif (CLK'event and CLK='1') then
      if (CLKEN='1') then 
			  IQ <= D;
		  end if;
    end if;
	 
    if OE = '1' then 
      if (CLK'event and CLK='0') then
		    Q <= IQ;
      end if;
    else
		  Q <= (others => 'Z');
	  end if;
	
  end process;
end arch;